module cobra (
  input clk,
  input up,
  input down,
  input left,
  input right,
  output [1:0] next_pos
);

endmodule
