module fruta #(
    parameter MAPA_HEIGHT,
    parameter MAPA_WIDTH
) (
    input [1:0] mapa_dado,
    output [9:0] mapa_x,
    output [9:0] mapa_y,
    output mapa_read,
    output mapa_write
);

    
endmodule //fruta